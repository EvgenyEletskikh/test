`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// �����������: ��� ����
// ��������: ������� ������� ���������
// ���������: ������� ������ ���-42
// 
// �������� �������: ���������� ��������� CORDIC ��� ���������� ���������� ����� ��������������� ����� � �������
// �������� ������: tb.v
//
// ������ ���������: Vivado 2019.1
// 
// ��������:
//      ������ ������� �� ���� ������:
//          1) ������ tb.v - �������� ��� ������������ ������ �������
//          2) ������ cordic_top.v - ������, ����������� �� ���� �������� � ����� ������ ��������� (���������� 
//                  ���������������� ������, ���������������� �������� ��� ����������) � ����������� 16-��� �������
//                  cordic-unit ��� ����������� ������������ ����������
//          3) ������ cordic_unit.v - ������, ����������� ������������� ��� � ���������, ��������������� �������������
//                  � �������� ��������� ������ �������� 
//////////////////////////////////////////////////////////////////////////////////

module tb();

reg CLK;
reg [7:0] loopy;

reg signed [31:0] ix,iy,iz;
wire signed [31:0] out;

parameter ITERS = 16;
parameter SW = 3;

cordic_top #(ITERS,SW) dut(
                    .CLK(CLK),
                    .ix(ix),
                    .iy(iy),     
                    .iz(iz),       
                    .Res(out)
                    );
    
integer iter;        
initial begin
    CLK = 0;
    loopy = 0;
    for (iter = 0; iter < 40; iter = iter+1) begin
        #1 CLK = ~CLK;
        #1 CLK = ~CLK;
        loopy = loopy + 1;
    end
    $finish;
end

initial begin
    ix = 0;
    iy = 0;
    /*
    #1.5 // sh(-1.00) = -1.08620123136814084042
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111110000000000000000; // z = -1.000000
    
    #2 // sh(-0.60) = -0.70699907196315636693
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111110110011001100110; // z = -0.600006
    
    #2 // sh(-0.20) = -0.26174320291462316312
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111111100110011001101; // z = -0.199997
    
    #2 // sh(0.20) = 0.26174320291462316312
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000000011001100110011; // z = 0.199997
    
    #2 // sh(0.60) = 0.70699907196315636693
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000001001100110011010; // z = 0.600006
    
    #2 // sh(1.00) = 1.08620123136814084042
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000010000000000000000; // z = 1.000000
    */
    /*
    #1.5 // ch(-1.00) = 1.47625458519979479988
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111110000000000000000; // z = -1.000000
    
    #2 // ch(-0.60) = 1.22447628521524154444
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111110110011001100110; // z = -0.600006
    
    #2 // ch(-0.20) = 1.03391700910631278987
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111111100110011001101; // z = -0.199997
    
    #2 // ch(0.20) = 1.03391700910631278987
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000000011001100110011; // z = 0.199997
    
    #2 // ch(0.60) = 1.22447628521524154444
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000001001100110011010; // z = 0.600006
    
    #2 // ch(1.00) = 1.47625458519979479988
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000010000000000000000; // z = 1.000000
    */
    
    #1.5 // exp(-1.00) = 0.39005335383165395946
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111110000000000000000; // z = -1.000000
    
    #2 // exp(-0.60) = 0.51747721325208517751
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111110110011001100110; // z = -0.600006
    
    #2 // exp(-0.20) = 0.77217380619168962674
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b11111111111111111100110011001101; // z = -0.199997
    
    #2 // exp(0.20) = 1.29566021202093595299
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000000011001100110011; // z = 0.199997
    
    #2 // exp(0.60) = 1.93147535717839780034
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000001001100110011010; // z = 0.600006
    
    #2 // exp(1.00) = 2.56245581656793586234
    ix = 32'b00000000000000010011010010000100; // x = 1.205139
    iy = 32'b0;
    iz = 32'b00000000000000010000000000000000; // z = 1.000000
    
    
    
    
    
    #2 // 25
    ix = 32'b0;
    iy = 32'b0;
    iz = 32'b0;
end


endmodule